module special(
    input [2:0]i, 
	 input [2:0]j, 
	 output [5:0]damage, 
	 output [2:0]move,
	 output [5:0]heal, 
	 output stun, 
	 output [2:0]cost);
	 
	 always @(*) begin
	  // grab memory
	 end
	 
endmodule 